module rvfi_wrapper (
	input         clock,
	input         reset,
	`RVFI_OUTPUTS
);


(* keep *) `rvformal_rand_reg [31:0] IMEM_rd_data_i;
(* keep *) `rvformal_rand_reg [31:0] DMEM_rd_data_i;
(* keep *) logic [31:0] IMEM_addr_o;
(* keep *) logic [31:0] DMEM_addr_o;
(* keep *) logic [31:0] DMEM_wr_data_o;
(* keep *) logic [3:0] DMEM_wr_byte_en_o;

    dtcore32  dtcore32_inst (
    .clk_i(clock),
    .rst_i(reset),
    .IMEM_rd_data_i(IMEM_rd_data_i),
    .DMEM_rd_data_i(DMEM_rd_data_i),
    .rvfi_valid(rvfi_valid),
    .rvfi_order(rvfi_order),
    .rvfi_insn(rvfi_insn),
    .rvfi_trap(rvfi_trap),
    .rvfi_halt(rvfi_halt),
    .rvfi_intr(rvfi_intr),
    .rvfi_mode(rvfi_mode),
    .rvfi_ixl(rvfi_ixl),
    .rvfi_rs1_addr(rvfi_rs1_addr),
    .rvfi_rs2_addr(rvfi_rs2_addr),
    .rvfi_rs1_rdata(rvfi_rs1_rdata),
    .rvfi_rs2_rdata(rvfi_rs2_rdata),
    .rvfi_rd_addr(rvfi_rd_addr),
    .rvfi_rd_wdata(rvfi_rd_wdata),
    .rvfi_pc_rdata(rvfi_pc_rdata),
    .rvfi_pc_wdata(rvfi_pc_wdata),
    .rvfi_mem_addr(rvfi_mem_addr),
    .rvfi_mem_rmask(rvfi_mem_rmask),
    .rvfi_mem_wmask(rvfi_mem_wmask),
    .rvfi_mem_rdata(rvfi_mem_rdata),
    .rvfi_mem_wdata(rvfi_mem_wdata),
    .rvfi_csr_mcycle_rmask(rvfi_csr_mcycle_rmask),
    .rvfi_csr_mcycle_wmask(rvfi_csr_mcycle_wmask),
    .rvfi_csr_mcycle_rdata(rvfi_csr_mcycle_rdata),
    .rvfi_csr_mcycle_wdata(rvfi_csr_mcycle_wdata),
    .rvfi_csr_minstret_rmask(rvfi_csr_minstret_rmask),
    .rvfi_csr_minstret_wmask(rvfi_csr_minstret_wmask),
    .rvfi_csr_minstret_rdata(rvfi_csr_minstret_rdata),
    .rvfi_csr_minstret_wdata(rvfi_csr_minstret_wdata),
    .IMEM_addr_o(IMEM_addr_o),
    .DMEM_addr_o(DMEM_addr_o),
    .DMEM_wr_data_o(DMEM_wr_data_o),
    .DMEM_wr_byte_en_o(DMEM_wr_byte_en_o)
  );
endmodule

