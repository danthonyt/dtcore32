//`define RISCV_FORMAL