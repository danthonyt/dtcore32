module trap_unit(
    
);
endmodule