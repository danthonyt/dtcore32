//===========================================================
// Project    : RISC-V CPU
// File       : regfile.sv
// Module     : regfile
// Description: CPU register file for general-purpose registers.
//              Supports two read ports and one write port, synchronous
//              writes, and asynchronous reads.
//
// Inputs:
//   clk_i           - System clock
//   rst_i           - Synchronous reset
//   write_en_i      - Write enable for destination register
//   rs1_addr_i      - Source register 1 address
//   rs2_addr_i      - Source register 2 address
//   rd_addr_i       - Destination register address
//   reg_wr_data_i   - Data to write into the destination register
//
// Outputs:
//   rs1_rdata_o     - Data read from source register 1
//   rs2_rdata_o     - Data read from source register 2
//
// Notes:
//   - Implements 32 general-purpose registers (x0–x31) for RISC-V.
//   - Register x0 is hardwired to zero and ignores writes.
//   - Asynchronous read allows combinational access to rs1_rdata_o and rs2_rdata_o.
//   - Fully synchronous write occurs on the rising edge of clk_i.
//
// Author     : David Torres
// Date       : 2025-09-16
//===========================================================

module regfile (
    input logic clk_i,
    input logic rst_i,

    input logic write_en_i,
    input  logic [ 4:0] rs1_addr_i,
    input  logic [ 4:0] rs2_addr_i,
    input  logic [ 4:0] rd_addr_i,
    input  logic [31:0] reg_wr_data_i,
    output logic [31:0] rs1_rdata_o,
    output logic [31:0] rs2_rdata_o
);
  integer i;
  logic [31:0] reg_array[0:31];

  // three ported register file
  // read two ports combinationally (A1/RD1, A2/RD2)
  // write third port on rising edge of clock (A3/WD3/WE3)
  // register 0 hardwired to 0
  always_ff @(posedge clk_i) begin
    if (rst_i) begin
      for (i = 0; i < 32; i = i + 1) reg_array[i] <= 32'd0;
    end else if (write_en_i)begin
      if (rd_addr_i != 0) reg_array[rd_addr_i] <= reg_wr_data_i;
    end
  end
    assign rs1_rdata_o = reg_array[rs1_addr_i];
    assign rs2_rdata_o = reg_array[rs2_addr_i];

endmodule

