module dtcore32_top (
    input  logic CLK,
    input  logic RST,
    input  logic RX,
    output logic TX

);
  logic rstn;
  assign rstn = ~RST;
  localparam WISHBONE_ADDR_WIDTH = 32;
  localparam WISHBONE_BUS_WIDTH = 32;

  reg [WISHBONE_ADDR_WIDTH-1:0] IMEM_CMD_ADDR_O;
  reg [ WISHBONE_BUS_WIDTH-1:0] IMEM_CMD_RDATA_I;
  reg MEM_CMD_START_O;
  reg MEM_CMD_WE_O;
  reg [WISHBONE_ADDR_WIDTH-1:0] MEM_CMD_ADDR_O;
  reg [WISHBONE_BUS_WIDTH-1:0] MEM_CMD_WDATA_O;
  reg [(WISHBONE_BUS_WIDTH/8)-1:0] MEM_CMD_SEL_O;
  reg [WISHBONE_BUS_WIDTH-1:0] MEM_CMD_RDATA_I;
  reg MEM_CMD_BUSY_I;



  dtcore32 # (
    .WISHBONE_ADDR_WIDTH(WISHBONE_ADDR_WIDTH),
    .WISHBONE_BUS_WIDTH(WISHBONE_BUS_WIDTH)
  )
  dtcore32_inst (
    .CLK(CLK),
    .RST(RST),
    .IMEM_CMD_ADDR_O(IMEM_CMD_ADDR_O),
    .IMEM_CMD_RDATA_I(IMEM_CMD_RDATA_I),
    .MEM_CMD_START_O(MEM_CMD_START_O),
    .MEM_CMD_WE_O(MEM_CMD_WE_O),
    .MEM_CMD_ADDR_O(MEM_CMD_ADDR_O),
    .MEM_CMD_WDATA_O(MEM_CMD_WDATA_O),
    .MEM_CMD_SEL_O(MEM_CMD_SEL_O),
    .MEM_CMD_RDATA_I(MEM_CMD_RDATA_I),
    .MEM_CMD_BUSY_I(MEM_CMD_BUSY_I)
  );
endmodule
