module trap_handler(

);
endmodule