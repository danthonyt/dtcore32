`define RISCV_FORMAL