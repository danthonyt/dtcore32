//===========================================================
// Project    : RISC-V CPU
// File       : dtcore32.v
// Module     : dtcore32
// Description: Top-level CPU core module implementing a 32-bit
//              RISC-V pipeline. Interfaces with instruction memory,
//              and a unified data interface for memory-mapped
//              data memory or peripherals. Handles CSR, traps, and
//              optional formal verification signals (`RISCV_FORMAL`).
//
// Inputs:
//   clk_i                - System clock
//   rst_i                - Synchronous reset
//   imem_rdata_i         - Instruction memory read data
//   mem_rdata_i          - Read data from data memory or peripheral
//   mem_done_i           - Transaction completion from data memory or peripheral
//   (RISCV_FORMAL) rvfi signals - Optional outputs for formal verification
//
// Outputs:
//   imem_addr_o          - Instruction memory address
//   mem_valid_o          - Valid signal for data memory or peripheral transaction
//   mem_wen_o            - Write enable for data memory or peripheral
//   mem_addr_o           - Address for data memory or peripheral
//   mem_wdata_o          - Write data for data memory or peripheral
//   mem_strb_o           - Byte-enable strobes for write operations
//   (RISCV_FORMAL) rvfi signals - Optional formal verification outputs
//
// Notes:
//   - Integrates instruction fetch, decode, execute, memory, and write-back stages.
//   - Unified `mem_*` interface can access both data memory and memory-mapped peripherals.
//   - Optional RISCV_FORMAL signals allow formal verification of CPU behavior.
//   - Designed to interface with external CSR module and trap handling logic.
//
// Author     : David Torres
// Date       : 2025-09-16
//===========================================================
import riscv_pkg::*;
// Optional: conditional compilation flag
`define RISCV_FORMAL
module dtcore32 (
  input             clk_i                  ,
  input             rst_i                  ,
`ifdef RISCV_FORMAL
  output reg        rvfi_valid             ,
  output reg [63:0] rvfi_order             ,
  output reg [31:0] rvfi_insn              ,
  output reg        rvfi_trap              ,
  output reg        rvfi_halt              ,
  output reg        rvfi_intr              ,
  output reg [ 1:0] rvfi_mode              ,
  output reg [ 1:0] rvfi_ixl               ,
  output reg [ 4:0] rvfi_rs1_addr          ,
  output reg [ 4:0] rvfi_rs2_addr          ,
  output reg [31:0] rvfi_rs1_rdata         ,
  output reg [31:0] rvfi_rs2_rdata         ,
  output reg [ 4:0] rvfi_rd_addr           ,
  output reg [31:0] rvfi_rd_wdata          ,
  output reg [31:0] rvfi_pc_rdata          ,
  output reg [31:0] rvfi_pc_wdata          ,
  output reg [31:0] rvfi_mem_addr          ,
  output reg [ 3:0] rvfi_mem_rmask         ,
  output reg [ 3:0] rvfi_mem_wmask         ,
  output reg [31:0] rvfi_mem_rdata         ,
  output reg [31:0] rvfi_mem_wdata         ,
  output reg [63:0] rvfi_csr_mcycle_rmask  ,
  output reg [63:0] rvfi_csr_mcycle_wmask  ,
  output reg [63:0] rvfi_csr_mcycle_rdata  ,
  output reg [63:0] rvfi_csr_mcycle_wdata  ,
  output reg [63:0] rvfi_csr_minstret_rmask,
  output reg [63:0] rvfi_csr_minstret_wmask,
  output reg [63:0] rvfi_csr_minstret_rdata,
  output reg [63:0] rvfi_csr_minstret_wdata,
  output reg [31:0] rvfi_csr_mcause_rmask  ,
  output reg [31:0] rvfi_csr_mcause_wmask  ,
  output reg [31:0] rvfi_csr_mcause_rdata  ,
  output reg [31:0] rvfi_csr_mcause_wdata  ,
  output reg [31:0] rvfi_csr_mepc_rmask    ,
  output reg [31:0] rvfi_csr_mepc_wmask    ,
  output reg [31:0] rvfi_csr_mepc_rdata    ,
  output reg [31:0] rvfi_csr_mepc_wdata    ,
  output reg [31:0] rvfi_csr_mtvec_rmask   ,
  output reg [31:0] rvfi_csr_mtvec_wmask   ,
  output reg [31:0] rvfi_csr_mtvec_rdata   ,
  output reg [31:0] rvfi_csr_mtvec_wdata   ,
`endif
  // to instruction memory interface
  input      [31:0] imem_rdata_i           ,
  output reg [31:0] imem_addr_o            ,
  // to data memory and peripheral interface
  input      [31:0] mem_rdata_i            ,
  input             mem_done_i             ,
  output            mem_valid_o            ,
  output reg        mem_wen_o              ,
  output reg [31:0] mem_addr_o             ,
  output reg [31:0] mem_wdata_o            ,
  output reg [ 3:0] mem_strb_o
);


// ---------------- IF/ID PIPELINE REGISTERS ----------------
// Going in / Coming out
  reg        if_d_valid, id_q_valid;
  reg [31:0] if_d_pc, id_q_pc;
  reg [31:0] if_d_pc_plus_4, id_q_pc_plus_4;
  reg [31:0] if_d_insn, id_q_insn;
`ifdef RISCV_FORMAL
  reg if_d_intr, id_q_intr;
`endif

// ---------------- ID/EX PIPELINE REGISTERS ----------------
// Going in / Coming out
  reg        id_d_valid, ex_q_valid;
  reg [31:0] id_d_pc, ex_q_pc;
  reg [31:0] id_d_pc_plus_4, ex_q_pc_plus_4;
  reg [ 4:0] id_d_rs1_addr, ex_q_rs1_addr;
  reg [ 4:0] id_d_rs2_addr, ex_q_rs2_addr;
  reg [ 4:0] id_d_rd_addr, ex_q_rd_addr;
  reg [31:0] id_d_rs1_rdata, ex_q_rs1_rdata;
  reg [31:0] id_d_rs2_rdata, ex_q_rs2_rdata;
  reg [31:0] id_d_imm_ext, ex_q_imm_ext;
  reg [11:0] id_d_csr_addr, ex_q_csr_addr;
  reg [31:0] id_d_csr_rdata, ex_q_csr_rdata;

  reg [       ALU_CTRL_T_WIDTH-1:0] id_d_alu_control, ex_q_alu_control;
  reg [      ALU_A_SEL_T_WIDTH-1:0] id_d_alu_a_sel, ex_q_alu_a_sel;
  reg [      ALU_B_SEL_T_WIDTH-1:0] id_d_alu_b_sel, ex_q_alu_b_sel;
  reg [     PC_ALU_SEL_T_WIDTH-1:0] id_d_pc_alu_sel, ex_q_pc_alu_sel;
  reg [CSR_BITMASK_SEL_T_WIDTH-1:0] id_d_csr_bitmask_sel, ex_q_csr_bitmask_sel;

  reg id_d_is_branch, ex_q_is_branch;
  reg id_d_is_jump, ex_q_is_jump;
  reg id_d_is_csr_write, ex_q_is_csr_write;
  reg id_d_is_csr_read, ex_q_is_csr_read;
  reg id_d_is_rd_write, ex_q_is_rd_write;
  reg id_d_is_rs1_read, ex_q_is_rs1_read;
  reg id_d_is_rs2_read, ex_q_is_rs2_read;
  reg id_d_is_mem_write, ex_q_is_mem_write;
  reg id_d_is_mem_read, ex_q_is_mem_read;

  reg id_d_is_jal, ex_q_is_jal;
  reg id_d_is_jalr, ex_q_is_jalr;
  reg id_d_is_memsize_b, ex_q_is_memsize_b;
  reg id_d_is_memsize_bu, ex_q_is_memsize_bu;
  reg id_d_is_memsize_h, ex_q_is_memsize_h;
  reg id_d_is_memsize_hu, ex_q_is_memsize_hu;
  reg id_d_is_memsize_w, ex_q_is_memsize_w;

  reg id_d_csr_op_rw, ex_q_csr_op_rw;
  reg id_d_csr_op_clear, ex_q_csr_op_clear;
  reg id_d_csr_op_set, ex_q_csr_op_set;

  reg       id_d_branch_predict, ex_q_branch_predict;
  reg [5:0] id_d_pht_idx, ex_q_pht_idx;

  reg        id_d_trap_valid, ex_q_trap_valid;
  reg [31:0] id_d_trap_mcause, ex_q_trap_mcause;
  reg [31:0] id_d_trap_pc, ex_q_trap_pc;

`ifdef RISCV_FORMAL
  reg [31:0] id_d_insn, ex_q_insn;
  reg        id_d_intr, ex_q_intr;
// For rvfi_trap_info, you can either flatten all fields or leave as separate regs
  reg [31:0] id_d_trap_insn,     ex_q_trap_insn;
  reg [31:0] id_d_trap_next_pc,  ex_q_trap_next_pc;
  reg [ 4:0] id_d_trap_rs1_addr, ex_q_trap_rs1_addr;
  reg [ 4:0] id_d_trap_rs2_addr, ex_q_trap_rs2_addr;
  reg [ 4:0] id_d_trap_rd_addr,  ex_q_trap_rd_addr;
  reg [31:0] id_d_trap_rs1_rdata, ex_q_trap_rs1_rdata;
  reg [31:0] id_d_trap_rs2_rdata, ex_q_trap_rs2_rdata;
  reg [31:0] id_d_trap_rd_wdata, ex_q_trap_rd_wdata;

`endif
// ---------------- EX/MEM PIPELINE REGISTERS ----------------
// Going in / Coming out
  reg        ex_d_valid,          mem_q_valid;
  reg [31:0] ex_d_pc,             mem_q_pc;
  reg [31:0] ex_d_pc_plus_4,      mem_q_pc_plus_4;
  reg [ 4:0] ex_d_rd_addr,        mem_q_rd_addr;
  reg [11:0] ex_d_csr_addr,       mem_q_csr_addr;
  reg [31:0] ex_d_csr_wdata,      mem_q_csr_wdata;

  reg [31:0] ex_d_store_wdata,    mem_q_store_wdata;
  reg [31:0] ex_d_alu_csr_result, mem_q_alu_csr_result;

  reg ex_d_is_branch,      mem_q_is_branch;
  reg ex_d_is_jump,        mem_q_is_jump;
  reg ex_d_is_csr_write,   mem_q_is_csr_write;
  reg ex_d_is_csr_read,    mem_q_is_csr_read;
  reg ex_d_is_rd_write,    mem_q_is_rd_write;
  reg ex_d_is_mem_write,   mem_q_is_mem_write;
  reg ex_d_is_mem_read,    mem_q_is_mem_read;

  reg ex_d_is_jal,         mem_q_is_jal;
  reg ex_d_is_jalr,        mem_q_is_jalr;
  reg ex_d_is_memsize_b,   mem_q_is_memsize_b;
  reg ex_d_is_memsize_bu,  mem_q_is_memsize_bu;
  reg ex_d_is_memsize_h,   mem_q_is_memsize_h;
  reg ex_d_is_memsize_hu,  mem_q_is_memsize_hu;
  reg ex_d_is_memsize_w,   mem_q_is_memsize_w;

  reg       ex_d_branch_predict, mem_q_branch_predict;
  reg [5:0] ex_d_pht_idx,        mem_q_pht_idx;

  reg        ex_d_jump_taken,     mem_q_jump_taken;
  reg [31:0] ex_d_jaddr,          mem_q_jaddr;

  reg        ex_d_trap_valid,     mem_q_trap_valid;
  reg [31:0] ex_d_trap_mcause,    mem_q_trap_mcause;
  reg [31:0] ex_d_trap_pc,        mem_q_trap_pc;

`ifdef RISCV_FORMAL
  reg [31:0] ex_d_insn,           mem_q_insn;
  reg        ex_d_intr,           mem_q_intr;
  reg [31:0] ex_d_next_pc,        mem_q_next_pc;
  reg [31:0] ex_d_csr_rdata,      mem_q_csr_rdata;
  reg [ 4:0] ex_d_rs1_addr,       mem_q_rs1_addr;
  reg [ 4:0] ex_d_rs2_addr,       mem_q_rs2_addr;
  reg [31:0] ex_d_rs1_rdata,      mem_q_rs1_rdata;
  reg [31:0] ex_d_rs2_rdata,      mem_q_rs2_rdata;
// Flattened trap_info_t inside ex_mem_t
  reg [31:0] ex_d_trap_insn,      mem_q_trap_insn;
  reg [31:0] ex_d_trap_next_pc,   mem_q_trap_next_pc;
  reg [ 4:0] ex_d_trap_rs1_addr,  mem_q_trap_rs1_addr;
  reg [ 4:0] ex_d_trap_rs2_addr,  mem_q_trap_rs2_addr;
  reg [ 4:0] ex_d_trap_rd_addr,   mem_q_trap_rd_addr;
  reg [31:0] ex_d_trap_rs1_rdata, mem_q_trap_rs1_rdata;
  reg [31:0] ex_d_trap_rs2_rdata, mem_q_trap_rs2_rdata;
  reg [31:0] ex_d_trap_rd_wdata,  mem_q_trap_rd_wdata;
`endif

// ---------------- MEM/WB PIPELINE REGISTERS ----------------
// Going in / Coming out
  reg        mem_d_valid,        wb_q_valid;
  reg [ 4:0] mem_d_rd_addr,      wb_q_rd_addr;
  reg [11:0] mem_d_csr_addr,     wb_q_csr_addr;
  reg [31:0] mem_d_csr_wdata,    wb_q_csr_wdata;
  reg [31:0] mem_d_rd_wdata,     wb_q_rd_wdata;
  reg [31:0] mem_d_pc_plus_4,    wb_q_pc_plus_4;

  reg mem_d_is_csr_write, wb_q_is_csr_write;
  reg mem_d_is_csr_read,  wb_q_is_csr_read;
  reg mem_d_is_rd_write,  wb_q_is_rd_write;

  reg        mem_d_trap_valid,   wb_q_trap_valid;
  reg [31:0] mem_d_trap_mcause,  wb_q_trap_mcause;
  reg [31:0] mem_d_trap_pc,      wb_q_trap_pc;

`ifdef RISCV_FORMAL
  reg [31:0] mem_d_pc,           wb_q_pc;
  reg [31:0] mem_d_next_pc,      wb_q_next_pc;
  reg [31:0] mem_d_insn,         wb_q_insn;
  reg        mem_d_intr,         wb_q_intr;
  reg [31:0] mem_d_csr_rdata,    wb_q_csr_rdata;
  reg [31:0] mem_d_mem_addr,     wb_q_mem_addr;
  reg [31:0] mem_d_load_rdata,   wb_q_load_rdata;
  reg [ 4:0] mem_d_rs1_addr,     wb_q_rs1_addr;
  reg [ 4:0] mem_d_rs2_addr,     wb_q_rs2_addr;
  reg [31:0] mem_d_rs1_rdata,    wb_q_rs1_rdata;
  reg [31:0] mem_d_rs2_rdata,    wb_q_rs2_rdata;
  reg [ 3:0] mem_d_load_rmask,   wb_q_load_rmask;
  reg [ 3:0] mem_d_store_wmask,  wb_q_store_wmask;
  reg [31:0] mem_d_store_wdata,  wb_q_store_wdata;
// Flattened trap_info_t inside mem_wb_t
  reg [31:0] mem_d_trap_insn,    wb_q_trap_insn;
  reg [31:0] mem_d_trap_next_pc, wb_q_trap_next_pc;
  reg [ 4:0] mem_d_trap_rs1_addr,wb_q_trap_rs1_addr;
  reg [ 4:0] mem_d_trap_rs2_addr,wb_q_trap_rs2_addr;
  reg [ 4:0] mem_d_trap_rd_addr, wb_q_trap_rd_addr;
  reg [31:0] mem_d_trap_rs1_rdata, wb_q_trap_rs1_rdata;
  reg [31:0] mem_d_trap_rs2_rdata, wb_q_trap_rs2_rdata;
  reg [31:0] mem_d_trap_rd_wdata, wb_q_trap_rd_wdata;
`endif


// ---------------- WB/RVFI PIPELINE REGISTERS ----------------
// Coming out



  wire if_id_stall;
  wire if_id_flush;

  wire id_ex_stall;
  wire id_ex_flush;

  wire ex_mem_stall;
  wire ex_mem_flush;

  wire mem_wb_stall;
  wire mem_wb_flush;
`ifdef RISCV_FORMAL

  wire [31:0] wb_csr_rmask;
  wire [31:0] wb_csr_wmask;
`endif
  // if stage signals;
  reg [31:0] next_pc          ;
  reg [31:0] trap_handler_addr;
  reg [31:0] imem_addr_q      ;
  reg        imem_rdata_valid ;
  reg        imem_buf_valid   ;
  reg [31:0] if_insn_buf      ;
  reg [31:0] if_buf_pc        ;
  // branch prediction logic
  wire [31:0] id_branch_addr   ;
  wire        id_predict_btaken;
  wire [ 5:0] id_pht_idx       ;
  // id stage signals
  wire                               id_forward_rs1       ;
  wire                               id_forward_rs2       ;
  reg  [                       11:0] id_csr_addr          ;
  reg  [                       31:0] id_imm_ext           ;
  reg  [                        4:0] id_rd_addr           ;
  wire [       ALU_CTRL_T_WIDTH-1:0] id_alu_control       ;
  reg  [                        6:0] id_op                ;
  reg  [                        2:0] id_funct3            ;
  reg                                id_funct7b5          ;
  reg  [                        6:0] id_funct7            ;
  reg  [                       11:0] id_funct12           ;
  reg                                id_rtype_alt         ;
  reg                                id_itype_alt         ;
  wire [     IMM_EXT_OP_T_WIDTH-1:0] id_imm_ext_op        ;
  wire [      ALU_A_SEL_T_WIDTH-1:0] id_alu_a_sel         ;
  wire [      ALU_B_SEL_T_WIDTH-1:0] id_alu_b_sel         ;
  wire [     PC_ALU_SEL_T_WIDTH-1:0] id_pc_alu_sel        ;
  wire [CSR_BITMASK_SEL_T_WIDTH-1:0] id_csr_bitmask_sel   ;
  reg  [                        4:0] id_rs1_addr          ;
  reg  [                        4:0] id_rs2_addr          ;
  wire [                       31:0] regfile_rs1_rdata    ;
  wire [                       31:0] regfile_rs2_rdata    ;
  reg  [                       31:0] csrfile_rdata        ;
  wire                               id_illegal_instr_trap;
  wire                               id_ecall_m_trap      ;
  wire                               id_breakpoint_trap   ;
  wire                               id_is_branch         ;
  wire                               id_is_jump           ;
  wire                               id_is_csr_write      ;
  wire                               id_is_csr_read       ;
  wire                               id_is_rd_write       ;
  wire                               id_is_rs1_read       ;
  wire                               id_is_rs2_read       ;
  wire                               id_is_mem_write      ;
  wire                               id_is_mem_read       ;
  wire                               id_is_jal            ;
  wire                               id_is_jalr           ;
  wire                               id_is_memsize_b      ;
  wire                               id_is_memsize_bu     ;
  wire                               id_is_memsize_h      ;
  wire                               id_is_memsize_hu     ;
  wire                               id_is_memsize_w      ;
  wire                               id_csr_op_rw         ;
  wire                               id_csr_op_clear      ;
  wire                               id_csr_op_set        ;

  // ex stage signal
  reg  [ 1:0] ex_forward_rs1_sel;
  reg  [ 1:0] ex_forward_rs2_sel;
  wire [31:0] ex_jaddr          ;
  wire        ex_jump_taken     ;
  reg  [31:0] ex_rs1_rdata      ;
  reg  [31:0] ex_rs2_rdata      ;
  reg  [31:0] ex_csr_bitmask    ;
  reg  [31:0] ex_csr_wdata      ;
  reg  [31:0] ex_src_a          ;
  reg  [31:0] ex_src_b          ;
  reg  [31:0] ex_pc_base        ;
  reg         ex_branch_cond    ;
  wire        ex_misaligned_jump;
  reg  [31:0] ex_alu_result     ;

  //mem stage
  reg         misaligned_load       ;
  reg         misaligned_store      ;
  reg  [ 3:0] mem_wstrb             ;
  reg  [ 3:0] mem_rstrb             ;
  reg         dmem_periph_req       ;
  reg  [31:0] mem_load_rdata        ;
  wire        mem_btaken_mispredict ;
  wire        mem_bntaken_mispredict;
  wire        mem_branch_mispredict ;
  // writeback stage
  reg [ 4:0] wb_rd_addr    ;
  reg [11:0] wb_csr_addr   ;
  reg [31:0] wb_rd_wdata   ;
  reg [31:0] wb_csr_wdata  ;
  reg [31:0] wb_trap_mcause;
  reg [31:0] wb_trap_pc    ;
  //*****************************************************************
  //
  //
  // INSTRUCTION FETCH STAGE
  //
  //
  //*****************************************************************

  // send read address to the instruction memory
  always @(posedge clk_i)
    begin
      if (rst_i)
        begin
          imem_addr_o      <= RESET_PC;
          imem_rdata_valid <= 0;
        end
      else if (if_id_flush) begin
        imem_addr_o      <= next_pc;
        imem_rdata_valid <= 0;
      end
      else if (!if_id_stall)
        begin
          imem_addr_o      <= next_pc;
          imem_rdata_valid <= 1;
        end
    end


  // registers imem address to stay cycle aligned with imem rdata
  // imem reads have 1 cycle latency
  always @(posedge clk_i)
    begin
      if (rst_i) begin
        imem_addr_q <= RESET_PC;
      end else begin
        imem_addr_q <= imem_addr_o;
      end
    end

  // buffer
  always @(posedge clk_i)
    begin
      if (rst_i)
        begin
          imem_buf_valid <= 0;
        end
      else if (if_id_flush) begin
        imem_buf_valid <= 0;
      end
      else if (!if_id_stall)
        begin
          imem_buf_valid <= 0;
        end
      // When entering a stall, buffer the instruction memory read data.
      // When first leaving a stall, use the buffered data instead. This
      // is to avoid losing instruction data when entering a stall.
      else if (if_id_stall && !imem_buf_valid)
        begin
          if_insn_buf    <= imem_rdata_i;
          imem_buf_valid <= 1;
          if_buf_pc      <= imem_addr_q;
        end
    end

  always @(*)
    begin
      // jump to trap handler if a trap instruction commits
      // else if a branch taken and mispredicted jump to mem.pc + 4
      // else if a branch not taken and mispredicted OR a jump instruction
      // jump to mem.jaddr
      // else if a branch taken is predicted jump to that address
      // else increment pc by 4
      next_pc = wb_q_trap_valid ? trap_handler_addr :
        mem_btaken_mispredict ? mem_q_pc_plus_4 :
        mem_bntaken_mispredict ? mem_q_jaddr :
        mem_q_jump_taken && !mem_q_is_branch ? mem_q_jaddr :
        id_predict_btaken ? id_branch_addr :
        imem_addr_o + 4;
      if_d_pc        = imem_buf_valid ? if_buf_pc : imem_addr_q;
      if_d_pc_plus_4 = if_d_pc + 4;
      if_d_insn      = imem_buf_valid ? if_insn_buf : imem_rdata_i;
      if_d_valid     = imem_rdata_valid;
    end

`ifdef RISCV_FORMAL
  reg if_intr_d ;
  reg if_intr_q ;
  reg if_intr_qq;
  always @(posedge clk_i)
    begin
      if (rst_i)
        begin
          if_intr_q  <= 0;
          if_intr_qq <= 0;
        end
      else if (if_id_flush)
        begin
          if_intr_q  <= 0;
          if_intr_qq <= 0;
        end
      else if (!if_id_stall)
        begin
          if_intr_q  <= if_intr_d;
          if_intr_qq <= if_intr_q;
        end
    end
  always @(*)
    begin
      if_d_intr = if_intr_qq;
      if_intr_d = wb_q_trap_valid;
    end
`endif
  //*****************************************************************
  //
  //
  // INSTRUCTION DECODE STAGE
  //
  //
  //*****************************************************************

  //*****************************************************************
  //
  //
  // GSHARE BRANCH PREDICTOR
  //
  //
  //*****************************************************************
  branch_predictor  branch_predictor_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .id_is_branch(id_is_branch),
    .id_q_pc(id_q_pc),
    .mem_q_is_branch(mem_q_is_branch),
    .mem_q_jump_taken(mem_q_jump_taken),
    .mem_q_pht_idx(mem_q_pht_idx),
    .id_predict_btaken(id_predict_btaken),
    .id_pht_idx(id_pht_idx)
  );

  reg illegal_instr_trap;
  reg ecall_m_trap      ;
  reg breakpoint_trap   ;

  reg is_branch    ;
  reg is_jump      ;
  reg is_jal       ;
  reg is_jalr      ;
  reg is_csr_write ;
  reg is_csr_read  ;
  reg csr_op_rw    ;
  reg csr_op_clear ;
  reg csr_op_set   ;
  reg is_rd_write  ;
  reg is_rs1_read  ;
  reg is_rs2_read  ;
  reg is_mem_write ;
  reg is_mem_read  ;
  reg is_memsize_b ;
  reg is_memsize_bu;
  reg is_memsize_h ;
  reg is_memsize_hu;
  reg is_memsize_w ;


  reg [       ALU_CTRL_T_WIDTH-1:0] alu_control    ;
  reg [     IMM_EXT_OP_T_WIDTH-1:0] imm_ext_op     ;
  reg [      ALU_A_SEL_T_WIDTH-1:0] alu_a_src      ;
  reg [      ALU_B_SEL_T_WIDTH-1:0] alu_b_src      ;
  reg [     PC_ALU_SEL_T_WIDTH-1:0] pc_alu_src     ;
  reg [CSR_BITMASK_SEL_T_WIDTH-1:0] csr_bitmask_sel;

  reg  [ALU_OP_T_WIDTH-1:0] alu_op                ;
  wire                      is_itype              ;
  wire                      is_rtype              ;
  wire                      is_SRAI_funct3        ;
  wire                      is_SRA_or_SUB_funct3  ;
  wire                      is_SLLI_or_SRLI_funct3;
  wire                      is_shift_itype        ;
  wire                      is_unknown_rtype      ;
  wire                      is_unknown_itype      ;

  assign is_itype               = (id_op == OPCODE_I_TYPE);
  assign is_rtype               = (id_op == OPCODE_R_TYPE);
  assign is_SRAI_funct3         = (id_funct3 == FUNCT3_SRAI);
  assign is_SRA_or_SUB_funct3   = ((id_funct3 == FUNCT3_SRA) || (id_funct3 == FUNCT3_SUB));
  assign is_SLLI_or_SRLI_funct3 = ((id_funct3 == FUNCT3_SLLI) || (id_funct3 == FUNCT3_SRLI));
  assign is_shift_itype         = is_SLLI_or_SRLI_funct3 | is_SRAI_funct3;
  assign is_unknown_rtype       = is_rtype
    & (id_funct7 != 7'h00)
    & ~((id_funct7 == 7'h20) & is_SRA_or_SUB_funct3);
  assign is_unknown_itype = is_itype
    & is_shift_itype
    & ~(is_SLLI_or_SRLI_funct3 & (id_funct7 == 7'h00))
    & ~(is_SRAI_funct3 & (id_funct7 == 7'h20));


  // Decode the control signals for the specific instruction
  always @(*) begin
    ecall_m_trap       = 0;
    illegal_instr_trap = 0;
    breakpoint_trap    = 0;
    // valid registers
    is_rd_write        = 0;
    is_rs1_read        = 0;
    is_rs2_read        = 0;
    // mux select signals
    alu_op             = 0;
    // control signals
    is_branch          = 0;
    is_jump            = 0;
    is_jal             = 0;
    is_jalr            = 0;
    is_csr_write       = 0;
    is_csr_read        = 0;
    csr_op_rw          = 0;
    csr_op_clear       = 0;
    csr_op_set         = 0;
    is_mem_write       = 0;
    is_mem_read        = 0;
    is_memsize_b       = 0;
    is_memsize_bu      = 0;
    is_memsize_h       = 0;
    is_memsize_hu      = 0;
    is_memsize_w       = 0;
    // sources
    imm_ext_op         = 0;
    alu_a_src          = 0;
    alu_b_src          = 0;
    pc_alu_src         = 0;
    csr_bitmask_sel    = 0;


    case (id_op)
      OPCODE_LOAD : begin
        imm_ext_op = I_ALU_TYPE;
        alu_a_src  = ALU_A_SEL_REG_DATA;
        alu_b_src  = ALU_B_SEL_IMM;
        alu_op     = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src = PC_ALU_SEL_PC;
        case (id_funct3)
          FUNCT3_LB : begin
            {is_rd_write, is_rs1_read, is_mem_read, is_memsize_b} = 4'b1111;
          end
          FUNCT3_LH : begin
            {is_rd_write, is_rs1_read, is_mem_read, is_memsize_h} = 4'b1111;
          end
          FUNCT3_LW : begin
            {is_rd_write, is_rs1_read, is_mem_read, is_memsize_w} = 4'b1111;
          end
          FUNCT3_LBU : begin
            {is_rd_write, is_rs1_read, is_mem_read, is_memsize_bu} = 4'b1111;
          end
          FUNCT3_LHU : begin
            {is_rd_write, is_rs1_read, is_mem_read, is_memsize_hu} = 4'b1111;
          end
          default : begin
            illegal_instr_trap = 1;
          end
        endcase
      end

      OPCODE_SYSCALL_CSR : begin
        case (id_funct3)
          FUNCT3_ECALL_EBREAK : begin
            if ((id_rs1_addr == 0) && (id_rd_addr == 0)) begin
              if (id_funct12 == 12'h001) begin
                breakpoint_trap = 1;
              end else if (id_funct12 == 12'h000) begin
                ecall_m_trap = 1;
              end else begin
                illegal_instr_trap = 1;
              end
            end else begin
              illegal_instr_trap = 1;
            end
          end
          // CSRRW/I always writes to the csr file, and conditionally reads when rd is not x0
          FUNCT3_CSRRW : begin
            {is_rs1_read, is_rd_write, is_csr_write, csr_op_rw} = 4'b1111;
            is_csr_read     = (id_rd_addr != 0);
            csr_bitmask_sel = CSR_BITMASK_SEL_REG_DATA;
          end
          FUNCT3_CSRRWI : begin
            {is_rs1_read, is_rd_write, is_csr_write, csr_op_rw} = 4'b1111;
            is_csr_read     = (id_rd_addr != 0);
            imm_ext_op      = CSR_TYPE;
            csr_bitmask_sel = CSR_BITMASK_SEL_IMM;
          end
          // Others always read from the csr file, and conditionally writes when
          // rs1 is x0, or uimm is 0 for register and immediate operand types, respectively
          FUNCT3_CSRRS : begin
            {is_rs1_read, is_rd_write, is_csr_read, csr_op_set} = 4'b1111;
            is_csr_write    = (id_rs1_addr != 0);
            csr_bitmask_sel = CSR_BITMASK_SEL_REG_DATA;
          end
          FUNCT3_CSRRSI : begin
            {is_rs1_read, is_rd_write, is_csr_read, csr_op_set} = 4'b1111;
            is_csr_write    = (id_rs1_addr != 0);
            imm_ext_op      = CSR_TYPE;
            csr_bitmask_sel = CSR_BITMASK_SEL_IMM;
          end
          FUNCT3_CSRRC : begin
            {is_rs1_read, is_rd_write, is_csr_read, csr_op_clear} = 4'b1111;
            is_csr_write    = (id_rs1_addr != 0);
            csr_bitmask_sel = CSR_BITMASK_SEL_REG_DATA;
          end
          FUNCT3_CSRRCI : begin
            {is_rs1_read, is_rd_write, is_csr_read, csr_op_clear} = 4'b1111;
            is_csr_write    = (id_rs1_addr != 0);
            imm_ext_op      = CSR_TYPE;
            csr_bitmask_sel = CSR_BITMASK_SEL_IMM;
          end
          default : begin
            illegal_instr_trap = 1;
          end
        endcase
      end
      OPCODE_STORE : begin
        imm_ext_op = S_TYPE;
        alu_a_src  = ALU_A_SEL_REG_DATA;
        alu_b_src  = ALU_B_SEL_IMM;
        alu_op     = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src = PC_ALU_SEL_PC;
        case (id_funct3)
          FUNCT3_SB : begin
            {is_rs1_read, is_rs2_read, is_mem_write, is_memsize_b} = 4'b1111;
          end
          FUNCT3_SH : begin
            {is_rs1_read, is_rs2_read, is_mem_write, is_memsize_h} = 4'b1111;
          end
          FUNCT3_SW : begin
            {is_rs1_read, is_rs2_read, is_mem_write, is_memsize_w} = 4'b1111;
          end
          default : begin
            illegal_instr_trap = 1;
          end
        endcase
      end
      OPCODE_R_TYPE : begin
        if (is_unknown_rtype) begin
          illegal_instr_trap = 1;
        end else begin
          {is_rs1_read, is_rs2_read, is_rd_write} = 3'b111;
          alu_a_src  = ALU_A_SEL_REG_DATA;
          alu_b_src  = ALU_B_SEL_REG_DATA;
          alu_op     = ALU_OP_IALU_ISHIFT_R_TYPE;
          pc_alu_src = PC_ALU_SEL_PC;
        end
      end
      OPCODE_B_TYPE : begin
        {is_rs1_read, is_rs2_read, is_branch} = 3'b111;
        imm_ext_op = B_TYPE;
        alu_a_src  = ALU_A_SEL_REG_DATA;
        alu_b_src  = ALU_B_SEL_REG_DATA;
        alu_op     = ALU_OP_B_TYPE;
        pc_alu_src = PC_ALU_SEL_PC;
      end
      //I-type ALU or shift
      OPCODE_I_TYPE : begin
        if (is_unknown_itype) begin
          illegal_instr_trap = 1;
        end else begin
          alu_a_src  = ALU_A_SEL_REG_DATA;
          alu_b_src  = ALU_B_SEL_IMM;
          alu_op     = ALU_OP_IALU_ISHIFT_R_TYPE;
          pc_alu_src = PC_ALU_SEL_PC;
          case (id_funct3)
            3'b000, 3'b010, 3'b011, 3'b100, 3'b110, 3'b111: begin
              {is_rs1_read, is_rd_write} = 2'b11;
              imm_ext_op = I_ALU_TYPE;  //I-type ALU
            end
            3'b001, 3'b101: begin
              {is_rs1_read, is_rd_write} = 2'b11;
              imm_ext_op = I_SHIFT_TYPE;  //I-type Shift
            end
            default : begin
              illegal_instr_trap = 1;
            end
          endcase  //I-type shift
        end
      end
      OPCODE_JAL : begin
        {is_rd_write, is_jump, is_jal} = 3'b111;
        imm_ext_op = J_TYPE;
        alu_a_src  = ALU_A_SEL_REG_DATA;
        alu_b_src  = ALU_B_SEL_REG_DATA;
        alu_op     = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src = PC_ALU_SEL_PC;
      end
      OPCODE_U_TYPE_LUI : begin
        is_rd_write = 1;
        imm_ext_op  = U_TYPE;
        alu_a_src   = ALU_A_SEL_ZERO;
        alu_b_src   = ALU_B_SEL_IMM;
        alu_op      = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src  = PC_ALU_SEL_PC;
      end
      OPCODE_U_TYPE_AUIPC : begin
        is_rd_write = 1;
        imm_ext_op  = U_TYPE;
        alu_a_src   = ALU_A_SEL_PC;
        alu_b_src   = ALU_B_SEL_IMM;
        alu_op      = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src  = PC_ALU_SEL_PC;
      end
      OPCODE_JALR : begin
        {is_rs1_read, is_rd_write, is_jump, is_jalr} = 4'b1111;
        imm_ext_op = I_ALU_TYPE;
        alu_a_src  = ALU_A_SEL_REG_DATA;
        alu_b_src  = ALU_B_SEL_IMM;
        alu_op     = ALU_OP_ILOAD_S_U_TYPE;
        pc_alu_src = PC_ALU_SEL_REG_DATA;
      end
      default : begin
        illegal_instr_trap = 1;
      end
    endcase
  end



  always @(*) begin
    alu_control = ADD_ALU_CONTROL;
    case (alu_op)
      //I-type Load, S-type, U-type
      ALU_OP_ILOAD_S_U_TYPE :
        alu_control = ADD_ALU_CONTROL;  //add- lw,sw,lb,lh,lbu,lhu,sb,sh,auipc,lui
      //B-type
      ALU_OP_B_TYPE :
        case (id_funct3)
          FUNCT3_BEQ  : alu_control = SUB_ALU_CONTROL;  //sub - beq
          FUNCT3_BNE  : alu_control = NE_ALU_CONTROL;  //sub - bne
          FUNCT3_BLT  : alu_control = LT_ALU_CONTROL;  //blt
          FUNCT3_BGE  : alu_control = GE_ALU_CONTROL;  //bge
          FUNCT3_BLTU : alu_control = LTU_ALU_CONTROL;  //bltu
          FUNCT3_BGEU : alu_control = GEU_ALU_CONTROL;  //bgeu
          default     : ;
        endcase
      //R-type, I-type ALU,I-type 1al shift
      ALU_OP_IALU_ISHIFT_R_TYPE : begin
        case (id_funct3)
          FUNCT3_ADD :
            alu_control = (id_rtype_alt) ? SUB_ALU_CONTROL  /*sub*/ : ADD_ALU_CONTROL  /*add*/;
          FUNCT3_SLL        : alu_control = L_SHIFT_ALU_CONTROL;  //sll
          FUNCT3_SLT        : alu_control = LT_ALU_CONTROL;  //slt
          FUNCT3_SLTU_SLTIU : alu_control = LTU_ALU_CONTROL;  //sltu, sltiu
          FUNCT3_XOR        : alu_control = XOR_ALU_CONTROL;  //xor
          FUNCT3_SRA        :
            alu_control = (id_rtype_alt || id_itype_alt) ? R_SHIFT_A_ALU_CONTROL /*sra*/ : R_SHIFT_L_ALU_CONTROL /*srl*/;
          FUNCT3_OR  : alu_control = OR_ALU_CONTROL;  //or
          FUNCT3_AND : alu_control = AND_ALU_CONTROL;  //and
          default    : ;
        endcase
      end
      default : ;
    endcase
  end

  assign id_alu_control        = alu_control;
  assign id_imm_ext_op         = imm_ext_op;
  assign id_alu_a_sel          = alu_a_src;
  assign id_alu_b_sel          = alu_b_src;
  assign id_pc_alu_sel         = pc_alu_src;
  assign id_csr_bitmask_sel    = csr_bitmask_sel;
  assign id_illegal_instr_trap = illegal_instr_trap;
  assign id_ecall_m_trap       = ecall_m_trap;
  assign id_breakpoint_trap    = breakpoint_trap;

  assign id_is_branch     = is_branch;
  assign id_is_jump       = is_jump;
  assign id_is_jal        = is_jal;
  assign id_is_jalr       = is_jalr;
  assign id_is_csr_write  = is_csr_write;
  assign id_is_csr_read   = is_csr_read;
  assign id_csr_op_rw     = csr_op_rw;
  assign id_csr_op_clear  = csr_op_clear;
  assign id_csr_op_set    = csr_op_set;
  assign id_is_rd_write   = (|id_rd_addr) ? is_rd_write : 0;
  assign id_is_rs1_read   = is_rs1_read;
  assign id_is_rs2_read   = is_rs2_read;
  assign id_is_mem_write  = is_mem_write;
  assign id_is_mem_read   = is_mem_read;
  assign id_is_memsize_b  = is_memsize_b;
  assign id_is_memsize_bu = is_memsize_bu;
  assign id_is_memsize_h  = is_memsize_h;
  assign id_is_memsize_hu = is_memsize_hu;
  assign id_is_memsize_w  = is_memsize_w;



riscv_imm_ext  riscv_imm_ext_inst (
    .id_q_insn(id_q_insn),
    .id_imm_ext_op(id_imm_ext_op),
    .id_imm_ext(id_imm_ext)
  );

  // compute branch address early to reduce combinational path of branch prediction
  assign id_branch_addr = id_q_pc +
    {{20{id_q_insn[31]}}, id_q_insn[7], id_q_insn[30:25], id_q_insn[11:8], 1'b0};
  // assign signals propagating to the next stage
  always @(*)
  begin
    id_op               = id_q_insn[6:0];
    id_funct3           = id_q_insn[14:12];
    id_funct7b5         = id_q_insn[30];
    id_funct7           = id_q_insn[31:25];
    id_funct12          = id_q_insn[31:20];
    id_rtype_alt        = id_op[5] & id_funct7b5;
    id_itype_alt        = ~id_op[5] & id_funct7b5;
    id_rs1_addr         = id_is_rs1_read ? id_q_insn[19:15] : 0;
    id_rs2_addr         = id_is_rs2_read ? id_q_insn[24:20] : 0;
    id_rd_addr          = id_q_insn[11:7];
    id_csr_addr         = id_q_insn[31:20];
    // Branch and jump
    id_d_is_branch      = id_is_branch;
    id_d_is_jump        = id_is_jump;
    id_d_is_jal         = id_is_jal;
    id_d_is_jalr        = id_is_jalr;
    id_d_branch_predict = id_predict_btaken;
    id_d_pht_idx        = id_pht_idx;

    // CSR operations
    id_d_is_csr_write = id_is_csr_write;
    id_d_is_csr_read  = id_is_csr_read;
    id_d_csr_op_rw    = id_csr_op_rw;
    id_d_csr_op_clear = id_csr_op_clear;
    id_d_csr_op_set   = id_csr_op_set;

    // Register reads/writes
    id_d_is_rd_write = id_is_rd_write;
    id_d_is_rs1_read = id_is_rs1_read;
    id_d_is_rs2_read = id_is_rs2_read;

    // Memory access
    id_d_is_mem_write = id_is_mem_write;
    id_d_is_mem_read  = id_is_mem_read;

    // Memory size indicators
    id_d_is_memsize_b  = id_is_memsize_b;
    id_d_is_memsize_bu = id_is_memsize_bu;
    id_d_is_memsize_h  = id_is_memsize_h;
    id_d_is_memsize_hu = id_is_memsize_hu;
    id_d_is_memsize_w  = id_is_memsize_w;

    //
    id_d_valid           = id_q_valid;
    id_d_pc              = id_q_pc;
    id_d_pc_plus_4       = id_q_pc_plus_4;
    id_d_rs1_addr        = id_rs1_addr;
    id_d_rs2_addr        = id_rs2_addr;
    id_d_rd_addr         = id_rd_addr;
    id_d_rs1_rdata       = id_forward_rs1 ? wb_rd_wdata : regfile_rs1_rdata;
    id_d_rs2_rdata       = id_forward_rs2 ? wb_rd_wdata : regfile_rs2_rdata;
    id_d_imm_ext         = id_imm_ext;
    id_d_csr_addr        = id_csr_addr;
    id_d_csr_rdata       = csrfile_rdata;
    id_d_alu_control     = id_alu_control;
    id_d_alu_a_sel       = id_alu_a_sel;
    id_d_alu_b_sel       = id_alu_b_sel;
    id_d_pc_alu_sel      = id_pc_alu_sel;
    id_d_csr_bitmask_sel = id_csr_bitmask_sel;
    // trap info
    if (id_ecall_m_trap) begin
      id_d_trap_valid  = 1;
      id_d_trap_pc     = id_q_pc;
      id_d_trap_mcause = {1'd0, TRAP_CODE_ECALL_M_MODE};
    end
    else if (id_breakpoint_trap) begin
      id_d_trap_valid  = 1;
      id_d_trap_pc     = id_q_pc;
      id_d_trap_mcause = {1'd0, TRAP_CODE_BREAKPOINT};
    end
    else if (id_illegal_instr_trap) begin
      id_d_trap_valid  = 1;
      id_d_trap_pc     = id_q_pc;
      id_d_trap_mcause = {1'd0, TRAP_CODE_ILLEGAL_INSTR};
    end
    else begin
      id_d_trap_valid  = 0;
      id_d_trap_mcause = 0;
      id_d_trap_pc     = 0;
    end

  end

`ifdef RISCV_FORMAL
  always @(*)
  begin
    // rvfi metadata
    id_d_insn           = id_q_insn;
    id_d_intr           = id_q_intr;
    // trap info for rvfi
    id_d_trap_insn      = id_q_insn;
    //id_d_trap_pc = id_q_pc;
    id_d_trap_next_pc   = 0;
    id_d_trap_rs1_addr  = 0;
    id_d_trap_rs2_addr  = 0;
    id_d_trap_rd_addr   = 0;
    id_d_trap_rs1_rdata = 0;
    id_d_trap_rs2_rdata = 0;
    id_d_trap_rd_wdata  = 0;
  end
`endif



  //*****************************************************************
  //
  //
  // INSTRUCTION EXECUTE STAGE
  //
  //
  //*****************************************************************

  // select rs1 read data
  always @(*) begin
    case (ex_forward_rs1_sel)
      NO_FORWARD_SEL :
        ex_rs1_rdata = ex_q_rs1_rdata;
      FORWARD_SEL_MEM_RESULT :
        ex_rs1_rdata = mem_q_alu_csr_result;
      FORWARD_SEL_WB_RESULT :
        ex_rs1_rdata = wb_rd_wdata;
      default :
        ex_rs1_rdata = 0;
    endcase
  end

// select input data for the first alu input
  always @(*) begin
    case (ex_q_alu_a_sel)
      ALU_A_SEL_REG_DATA :
        ex_src_a = ex_rs1_rdata;
      ALU_A_SEL_PC :
        ex_src_a = ex_q_pc;
      ALU_A_SEL_ZERO :
        ex_src_a = 0;
      default :
        ex_src_a = 0;
    endcase
  end

// select rs2 read data
  always @(*) begin
    case (ex_forward_rs2_sel)
      NO_FORWARD_SEL :
        ex_rs2_rdata = ex_q_rs2_rdata;
      FORWARD_SEL_MEM_RESULT :
        ex_rs2_rdata = mem_q_alu_csr_result;
      FORWARD_SEL_WB_RESULT :
        ex_rs2_rdata = wb_rd_wdata;
      default :
        ex_rs2_rdata = 0;
    endcase
  end

// select input data for the second alu input
  always @(*) begin
    case (ex_q_alu_b_sel)
      ALU_B_SEL_REG_DATA :
        ex_src_b = ex_rs2_rdata;
      ALU_B_SEL_IMM :
        ex_src_b = ex_q_imm_ext;
      default :
        ex_src_b = 0;
    endcase
  end

// select base value for pc offset
  always @(*) begin
    case (ex_q_pc_alu_sel)
      PC_ALU_SEL_REG_DATA :
        ex_pc_base = ex_rs1_rdata;
      PC_ALU_SEL_PC :
        ex_pc_base = ex_q_pc;
      default :
        ex_pc_base = 0;
    endcase
  end

// select bitmask source for csr op
  always @(*) begin
    case (ex_q_csr_bitmask_sel)
      CSR_BITMASK_SEL_REG_DATA :
        ex_csr_bitmask = ex_rs1_rdata;
      CSR_BITMASK_SEL_IMM :
        ex_csr_bitmask = ex_q_imm_ext;
      default :
        ex_csr_bitmask = 0;
    endcase
  end

// select csr result depending on op type
  always @(*) begin
    if (ex_q_csr_op_rw) begin
      ex_csr_wdata = ex_csr_bitmask;
    end
    else if (ex_q_csr_op_clear) begin
      ex_csr_wdata = (ex_q_csr_rdata & ~ex_csr_bitmask);
    end
    else if (ex_q_csr_op_set) begin
      ex_csr_wdata = (ex_q_csr_rdata | ex_csr_bitmask);
    end
    else begin
      ex_csr_wdata = 0;
    end
  end
  // trap if the jump address is not word aligned
  // jump if instruction is a jump or a branch and condition is true
  // jump is delayed to the mem stage to avoid long combinational path
  assign ex_jaddr           = (ex_q_is_jalr) ? ((ex_pc_base + ex_q_imm_ext) & ~(1'b1)) : (ex_pc_base + ex_q_imm_ext);
  assign ex_jump_taken      = (ex_q_is_jump | (ex_q_is_branch & ex_branch_cond));
  assign ex_misaligned_jump = ex_jump_taken & (ex_jaddr[1] | ex_jaddr[0]);

  always @(*)
    begin
      // Branch and jump
      ex_d_is_branch      = ex_q_is_branch;
      ex_d_is_jump        = ex_q_is_jump;
      ex_d_is_jal         = ex_q_is_jal;
      ex_d_is_jalr        = ex_q_is_jalr;
      ex_d_branch_predict = ex_q_branch_predict;
      ex_d_pht_idx        = ex_q_pht_idx;

      // CSR operations
      ex_d_is_csr_write = ex_q_is_csr_write;
      ex_d_is_csr_read  = ex_q_is_csr_read;

      // Register writes
      if (ex_misaligned_jump)
        ex_d_is_rd_write = 0;
      else
        ex_d_is_rd_write = ex_q_is_rd_write;

      // Memory access
      ex_d_is_mem_write = ex_q_is_mem_write;
      ex_d_is_mem_read  = ex_q_is_mem_read;

      // Memory size indicators
      ex_d_is_memsize_b  = ex_q_is_memsize_b;
      ex_d_is_memsize_bu = ex_q_is_memsize_bu;
      ex_d_is_memsize_h  = ex_q_is_memsize_h;
      ex_d_is_memsize_hu = ex_q_is_memsize_hu;
      ex_d_is_memsize_w  = ex_q_is_memsize_w;

      // pipeline
      ex_d_valid          = ex_q_valid;
      ex_d_pc             = ex_q_pc;
      ex_d_pc_plus_4      = ex_q_pc_plus_4;
      ex_d_rd_addr        = ex_q_rd_addr;
      ex_d_csr_addr       = ex_q_csr_addr;
      ex_d_csr_wdata      = ex_csr_wdata;
      ex_d_store_wdata    = ex_rs2_rdata;
      ex_d_alu_csr_result = (ex_q_is_csr_read) ? ex_q_csr_rdata : ex_alu_result;
      ex_d_jaddr          = ex_jaddr;
      ex_d_jump_taken     = ex_jump_taken;
      // traps
      if (ex_q_trap_valid)
        begin
          ex_d_trap_valid  = 1;
          ex_d_trap_mcause = ex_q_trap_mcause;
          ex_d_trap_pc     = ex_q_trap_pc;
        end
      else if (ex_misaligned_jump)
        begin
          ex_d_trap_valid  = 1;
          ex_d_trap_mcause = {1'b0, TRAP_CODE_INSTR_ADDR_MISALIGNED};
          ex_d_trap_pc     = ex_q_pc;
        end
      else
        begin
          ex_d_trap_valid  = 0;
          ex_d_trap_mcause = 0;
          ex_d_trap_pc     = 0;
        end
    end

  // calculates the branch condition of the instruction
  always @(*) begin
    case (ex_q_alu_control)
      SUB_ALU_CONTROL : ex_branch_cond = (ex_src_a == ex_src_b);  // beq
      NE_ALU_CONTROL  : ex_branch_cond = (ex_src_a != ex_src_b);
      LT_ALU_CONTROL  : ex_branch_cond = ($signed(ex_src_a) < $signed(ex_src_b));
      LTU_ALU_CONTROL : ex_branch_cond = (ex_src_a < ex_src_b);
      GE_ALU_CONTROL  : ex_branch_cond = ($signed(ex_src_a) >= $signed(ex_src_b));
      GEU_ALU_CONTROL : ex_branch_cond = (ex_src_a >= ex_src_b);
      default         : ex_branch_cond = 0;
    endcase
  end

  // calculates the result of the instruction
  always @(*) begin
    case (ex_q_alu_control)
      ADD_ALU_CONTROL       : ex_alu_result = ex_src_a + ex_src_b;
      SUB_ALU_CONTROL       : ex_alu_result = ex_src_a - ex_src_b;
      AND_ALU_CONTROL       : ex_alu_result = ex_src_a & ex_src_b;
      OR_ALU_CONTROL        : ex_alu_result = ex_src_a | ex_src_b;
      XOR_ALU_CONTROL       : ex_alu_result = ex_src_a ^ ex_src_b;
      LT_ALU_CONTROL, LTU_ALU_CONTROL: ex_alu_result = {31'd0, ex_branch_cond};
      L_SHIFT_ALU_CONTROL   : ex_alu_result = ex_src_a << ex_src_b[4:0];
      R_SHIFT_L_ALU_CONTROL : ex_alu_result = ex_src_a >> ex_src_b[4:0];
      R_SHIFT_A_ALU_CONTROL : ex_alu_result = $signed(ex_src_a) >>> ex_src_b[4:0];
      default               : ex_alu_result = 0;
    endcase
  end

`ifdef RISCV_FORMAL

  wire [31:0] ex_next_pc;
  assign ex_next_pc = (ex_jump_taken) ? ex_jaddr : ex_q_pc_plus_4;
  always @(*)
  begin
    // additional stage info
    ex_d_next_pc   = ex_next_pc;
    ex_d_insn      = ex_q_insn;
    ex_d_intr      = ex_q_intr;
    ex_d_rs1_addr  = ex_q_rs1_addr;
    ex_d_rs2_addr  = ex_q_rs2_addr;
    ex_d_rs1_rdata = ex_rs1_rdata;
    ex_d_rs2_rdata = ex_rs2_rdata;
    ex_d_csr_rdata = ex_q_csr_rdata;
    if (ex_q_trap_valid) // if trap from previous stage save it instead
      begin
        ex_d_trap_insn      = ex_q_trap_insn;
        ex_d_trap_next_pc   = ex_q_trap_next_pc;
        ex_d_trap_rs1_addr  = ex_q_trap_rs1_addr;
        ex_d_trap_rs2_addr  = ex_q_trap_rs2_addr;
        ex_d_trap_rd_addr   = ex_q_trap_rd_addr;
        ex_d_trap_rs1_rdata = ex_q_trap_rs1_rdata;
        ex_d_trap_rs2_rdata = ex_q_trap_rs2_rdata;
        ex_d_trap_rd_wdata  = ex_q_trap_rd_wdata;
      end else begin
      ex_d_trap_insn      = ex_q_insn;
      ex_d_trap_next_pc   = ex_next_pc;
      ex_d_trap_rs1_addr  = ex_q_rs1_addr;
      ex_d_trap_rs2_addr  = ex_q_rs2_addr;
      ex_d_trap_rd_addr   = ex_q_rd_addr;
      ex_d_trap_rs1_rdata = ex_src_a;
      ex_d_trap_rs2_rdata = ex_rs2_rdata;
      ex_d_trap_rd_wdata  = 0;
    end

  end
`endif
  //*****************************************************************
  //
  //
  // DATA MEMORY STAGE
  //
  //
  //*****************************************************************
  wire [4:0] load_size_onehot ;
  wire [2:0] store_size_onehot;
  wire       mem_valid        ;
  assign mem_btaken_mispredict  = (mem_q_is_branch && !mem_q_jump_taken && mem_q_branch_predict);
  assign mem_bntaken_mispredict = (mem_q_is_branch && mem_q_jump_taken && !mem_q_branch_predict);
  assign mem_branch_mispredict  = mem_btaken_mispredict || mem_bntaken_mispredict;
  assign load_size_onehot       = !mem_q_is_mem_read ? 0 :
    {
      mem_q_is_memsize_w,
      mem_q_is_memsize_hu,
      mem_q_is_memsize_h,
      mem_q_is_memsize_bu,
      mem_q_is_memsize_b
    };
  assign store_size_onehot = !mem_q_is_mem_write ? 0 :
    {
      mem_q_is_memsize_w,
      mem_q_is_memsize_h,
      mem_q_is_memsize_b
    };

  pulse_generator pulse_generator_inst (
    .clk_i  (clk_i                         ),
    .rst_i  (rst_i                         ),
    .en_i   (dmem_periph_req && !mem_done_i),
    .pulse_o(mem_valid                     )
  );
  assign mem_valid_o = mem_valid;
  //*****************************************************************
  //
  //
  // LOAD UNIT
  //
  //
  //*****************************************************************

load_unit  load_unit_inst (
    .mem_rdata_i(mem_rdata_i),
    .mem_q_alu_csr_result(mem_q_alu_csr_result),
    .load_size_onehot(load_size_onehot),
    .mem_rstrb(mem_rstrb),
    .mem_load_rdata(mem_load_rdata),
    .misaligned_load(misaligned_load)
  );

  //*****************************************************************
  //
  //
  // STORE UNIT
  //
  //
  //*****************************************************************
  store_unit  store_unit_inst (
    .mem_q_alu_csr_result(mem_q_alu_csr_result),
    .mem_q_store_wdata(mem_q_store_wdata),
    .store_size_onehot(store_size_onehot),
    .mem_wdata_o(mem_wdata_o),
    .mem_wstrb(mem_wstrb),
    .misaligned_store(misaligned_store)
  );

  always @(*)
    begin
      // memory interface local signals
      dmem_periph_req = (mem_q_is_mem_write || mem_q_is_mem_read) && !(misaligned_load || misaligned_store);
      mem_wen_o       = mem_q_is_mem_write;
      mem_addr_o      = mem_q_alu_csr_result;
      mem_strb_o      = mem_wen_o ? mem_wstrb : mem_rstrb;

      // pipeline
      mem_d_valid        = mem_q_valid;
      mem_d_is_csr_write = mem_q_is_csr_write;
      mem_d_is_csr_read  = mem_q_is_csr_read;
      mem_d_is_rd_write  = misaligned_load ? 0 : mem_q_is_rd_write;
      mem_d_rd_addr      = mem_q_rd_addr;
      mem_d_pc_plus_4    = mem_q_pc_plus_4;

      if (mem_q_is_jalr | mem_q_is_jal)  // is a jal or jalr
        mem_d_rd_wdata = mem_q_pc_plus_4;
      else if (mem_q_is_mem_read)  // is a load instruction
        mem_d_rd_wdata = mem_load_rdata;
      else  // else
        mem_d_rd_wdata = mem_q_alu_csr_result;

      mem_d_csr_addr  = mem_q_csr_addr;
      mem_d_csr_wdata = mem_q_csr_wdata;
      // traps
      if (mem_q_trap_valid)
        begin
          mem_d_trap_valid  = 1;
          mem_d_trap_mcause = mem_q_trap_mcause;
          mem_d_trap_pc     = mem_q_trap_pc;
        end
      else if (misaligned_store)
        begin
          mem_d_trap_valid  = 1;
          mem_d_trap_mcause = {1'b0, TRAP_CODE_STORE_ADDR_MISALIGNED};
          mem_d_trap_pc     = mem_q_pc;

        end
      else if (misaligned_load)
        begin
          mem_d_trap_valid  = 1;
          mem_d_trap_mcause = {1'b0, TRAP_CODE_LOAD_ADDR_MISALIGNED};
          mem_d_trap_pc     = mem_q_pc;
        end
      else
        begin
          mem_d_trap_valid  = 0;
          mem_d_trap_mcause = 0;
          mem_d_trap_pc     = 0;
        end
    end

`ifdef RISCV_FORMAL
  always @(*)
  begin
    // rvfi
    mem_d_pc      = mem_q_pc;
    // next pc changes on a branch mispredict
    mem_d_next_pc = mem_q_trap_valid ? trap_handler_addr :
      mem_q_jump_taken ? mem_q_jaddr :
      mem_q_pc_plus_4;
    mem_d_insn        = mem_q_insn;
    mem_d_intr        = mem_q_intr;
    mem_d_rs1_addr    = mem_q_rs1_addr;
    mem_d_rs2_addr    = mem_q_rs2_addr;
    mem_d_rs1_rdata   = mem_q_rs1_rdata;
    mem_d_rs2_rdata   = mem_q_rs2_rdata;
    // mem addresses are always word aligned
    mem_d_mem_addr    = mem_addr_o & ~32'h3;
    mem_d_load_rmask  = mem_rstrb;
    mem_d_store_wmask = mem_wstrb;
    mem_d_store_wdata = mem_wdata_o;
    mem_d_csr_rdata   = mem_q_csr_rdata;
    mem_d_load_rdata  = mem_rdata_i;
    // trap
    // if trap comes from previous stage save it instead
    if (mem_q_trap_valid) begin
      mem_d_trap_insn      = mem_q_trap_insn;
      mem_d_trap_next_pc   = mem_q_trap_next_pc;
      mem_d_trap_rs1_addr  = mem_q_trap_rs1_addr;
      mem_d_trap_rs2_addr  = mem_q_trap_rs2_addr;
      mem_d_trap_rd_addr   = mem_q_trap_rd_addr;
      mem_d_trap_rs1_rdata = mem_q_trap_rs1_rdata;
      mem_d_trap_rs2_rdata = mem_q_trap_rs2_rdata;
      mem_d_trap_rd_wdata  = 0;
    end else begin
      mem_d_trap_insn      = mem_q_insn;
      mem_d_trap_next_pc   = mem_q_next_pc;
      mem_d_trap_rs1_addr  = mem_q_rs1_addr;
      mem_d_trap_rs2_addr  = mem_q_rs2_addr;
      mem_d_trap_rd_addr   = mem_q_rd_addr;
      mem_d_trap_rs1_rdata = mem_q_rs1_rdata;
      mem_d_trap_rs2_rdata = mem_q_rs2_rdata;
      mem_d_trap_rd_wdata  = 0;
    end

  end
`endif

  //*****************************************************************
  //
  //
  // WRITEBACK STAGE
  //
  //
  //*****************************************************************


  always @(*)
    begin
      wb_trap_mcause = wb_q_trap_mcause;
      wb_trap_pc     = wb_q_trap_pc;
      wb_rd_addr     = wb_q_rd_addr;
      wb_rd_wdata    = wb_q_rd_wdata;
      wb_csr_addr    = wb_q_csr_addr;
      wb_csr_wdata   = wb_q_csr_wdata;
    end

  //*****************************************************************
  //
  //
  // PIPELINE REGISTERS
  //
  //
  //*****************************************************************


//-------------------------------
// IF/ID pipeline
//-------------------------------
if_id_pipeline  if_id_pipeline_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .if_id_flush(if_id_flush),
    .if_id_stall(if_id_stall),
    .imem_rdata_valid(imem_rdata_valid),
    .if_d_valid(if_d_valid),
    .if_d_pc(if_d_pc),
    .if_d_pc_plus_4(if_d_pc_plus_4),
    .if_d_insn(if_d_insn),
    .if_d_intr(if_d_intr),
    .id_q_intr(id_q_intr),
    .id_q_valid(id_q_valid),
    .id_q_pc(id_q_pc),
    .id_q_pc_plus_4(id_q_pc_plus_4),
    .id_q_insn(id_q_insn)
  );


//-------------------------------
// ID/EX pipeline
//-------------------------------
  id_ex_pipeline  id_ex_pipeline_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .id_ex_flush(id_ex_flush),
    .id_ex_stall(id_ex_stall),
    .if_id_stall(if_id_stall),
    .id_d_valid(id_d_valid),
    .id_d_pc(id_d_pc),
    .id_d_pc_plus_4(id_d_pc_plus_4),
    .id_d_rs1_addr(id_d_rs1_addr),
    .id_d_rs2_addr(id_d_rs2_addr),
    .id_d_rd_addr(id_d_rd_addr),
    .id_d_rs1_rdata(id_d_rs1_rdata),
    .id_d_rs2_rdata(id_d_rs2_rdata),
    .id_d_imm_ext(id_d_imm_ext),
    .id_d_csr_addr(id_d_csr_addr),
    .id_d_csr_rdata(id_d_csr_rdata),
    .id_d_alu_control(id_d_alu_control),
    .id_d_alu_a_sel(id_d_alu_a_sel),
    .id_d_alu_b_sel(id_d_alu_b_sel),
    .id_d_pc_alu_sel(id_d_pc_alu_sel),
    .id_d_csr_bitmask_sel(id_d_csr_bitmask_sel),
    .id_d_is_branch(id_d_is_branch),
    .id_d_is_jump(id_d_is_jump),
    .id_d_is_csr_write(id_d_is_csr_write),
    .id_d_is_csr_read(id_d_is_csr_read),
    .id_d_is_rd_write(id_d_is_rd_write),
    .id_d_is_rs1_read(id_d_is_rs1_read),
    .id_d_is_rs2_read(id_d_is_rs2_read),
    .id_d_is_mem_write(id_d_is_mem_write),
    .id_d_is_mem_read(id_d_is_mem_read),
    .id_d_is_jal(id_d_is_jal),
    .id_d_is_jalr(id_d_is_jalr),
    .id_d_is_memsize_b(id_d_is_memsize_b),
    .id_d_is_memsize_bu(id_d_is_memsize_bu),
    .id_d_is_memsize_h(id_d_is_memsize_h),
    .id_d_is_memsize_hu(id_d_is_memsize_hu),
    .id_d_is_memsize_w(id_d_is_memsize_w),
    .id_d_csr_op_rw(id_d_csr_op_rw),
    .id_d_csr_op_clear(id_d_csr_op_clear),
    .id_d_csr_op_set(id_d_csr_op_set),
    .id_d_branch_predict(id_d_branch_predict),
    .id_d_pht_idx(id_d_pht_idx),
    .id_d_trap_valid(id_d_trap_valid),
    .id_d_trap_mcause(id_d_trap_mcause),
    .id_d_trap_pc(id_d_trap_pc),
    .id_d_insn(id_d_insn),
    .id_d_intr(id_d_intr),
    .id_d_trap_insn(id_d_trap_insn),
    .id_d_trap_next_pc(id_d_trap_next_pc),
    .id_d_trap_rs1_addr(id_d_trap_rs1_addr),
    .id_d_trap_rs2_addr(id_d_trap_rs2_addr),
    .id_d_trap_rd_addr(id_d_trap_rd_addr),
    .id_d_trap_rs1_rdata(id_d_trap_rs1_rdata),
    .id_d_trap_rs2_rdata(id_d_trap_rs2_rdata),
    .id_d_trap_rd_wdata(id_d_trap_rd_wdata),
    .ex_q_insn(ex_q_insn),
    .ex_q_intr(ex_q_intr),
    .ex_q_trap_insn(ex_q_trap_insn),
    .ex_q_trap_next_pc(ex_q_trap_next_pc),
    .ex_q_trap_rs1_addr(ex_q_trap_rs1_addr),
    .ex_q_trap_rs2_addr(ex_q_trap_rs2_addr),
    .ex_q_trap_rd_addr(ex_q_trap_rd_addr),
    .ex_q_trap_rs1_rdata(ex_q_trap_rs1_rdata),
    .ex_q_trap_rs2_rdata(ex_q_trap_rs2_rdata),
    .ex_q_trap_rd_wdata(ex_q_trap_rd_wdata),
    .ex_q_valid(ex_q_valid),
    .ex_q_pc(ex_q_pc),
    .ex_q_pc_plus_4(ex_q_pc_plus_4),
    .ex_q_rs1_addr(ex_q_rs1_addr),
    .ex_q_rs2_addr(ex_q_rs2_addr),
    .ex_q_rd_addr(ex_q_rd_addr),
    .ex_q_rs1_rdata(ex_q_rs1_rdata),
    .ex_q_rs2_rdata(ex_q_rs2_rdata),
    .ex_q_imm_ext(ex_q_imm_ext),
    .ex_q_csr_addr(ex_q_csr_addr),
    .ex_q_csr_rdata(ex_q_csr_rdata),
    .ex_q_alu_control(ex_q_alu_control),
    .ex_q_alu_a_sel(ex_q_alu_a_sel),
    .ex_q_alu_b_sel(ex_q_alu_b_sel),
    .ex_q_pc_alu_sel(ex_q_pc_alu_sel),
    .ex_q_csr_bitmask_sel(ex_q_csr_bitmask_sel),
    .ex_q_is_branch(ex_q_is_branch),
    .ex_q_is_jump(ex_q_is_jump),
    .ex_q_is_csr_write(ex_q_is_csr_write),
    .ex_q_is_csr_read(ex_q_is_csr_read),
    .ex_q_is_rd_write(ex_q_is_rd_write),
    .ex_q_is_rs1_read(ex_q_is_rs1_read),
    .ex_q_is_rs2_read(ex_q_is_rs2_read),
    .ex_q_is_mem_write(ex_q_is_mem_write),
    .ex_q_is_mem_read(ex_q_is_mem_read),
    .ex_q_is_jal(ex_q_is_jal),
    .ex_q_is_jalr(ex_q_is_jalr),
    .ex_q_is_memsize_b(ex_q_is_memsize_b),
    .ex_q_is_memsize_bu(ex_q_is_memsize_bu),
    .ex_q_is_memsize_h(ex_q_is_memsize_h),
    .ex_q_is_memsize_hu(ex_q_is_memsize_hu),
    .ex_q_is_memsize_w(ex_q_is_memsize_w),
    .ex_q_csr_op_rw(ex_q_csr_op_rw),
    .ex_q_csr_op_clear(ex_q_csr_op_clear),
    .ex_q_csr_op_set(ex_q_csr_op_set),
    .ex_q_branch_predict(ex_q_branch_predict),
    .ex_q_pht_idx(ex_q_pht_idx),
    .ex_q_trap_valid(ex_q_trap_valid),
    .ex_q_trap_mcause(ex_q_trap_mcause),
    .ex_q_trap_pc(ex_q_trap_pc)
  );



//-------------------------------
// EX/MEM pipeline
//-------------------------------
  ex_mem_pipeline  ex_mem_pipeline_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .ex_mem_flush(ex_mem_flush),
    .ex_mem_stall(ex_mem_stall),
    .id_ex_stall(id_ex_stall),
    .ex_d_valid(ex_d_valid),
    .ex_d_pc(ex_d_pc),
    .ex_d_pc_plus_4(ex_d_pc_plus_4),
    .ex_d_rd_addr(ex_d_rd_addr),
    .ex_d_csr_addr(ex_d_csr_addr),
    .ex_d_csr_wdata(ex_d_csr_wdata),
    .ex_d_store_wdata(ex_d_store_wdata),
    .ex_d_alu_csr_result(ex_d_alu_csr_result),
    .ex_d_is_branch(ex_d_is_branch),
    .ex_d_is_jump(ex_d_is_jump),
    .ex_d_is_csr_write(ex_d_is_csr_write),
    .ex_d_is_csr_read(ex_d_is_csr_read),
    .ex_d_is_rd_write(ex_d_is_rd_write),
    .ex_d_is_mem_write(ex_d_is_mem_write),
    .ex_d_is_mem_read(ex_d_is_mem_read),
    .ex_d_is_jal(ex_d_is_jal),
    .ex_d_is_jalr(ex_d_is_jalr),
    .ex_d_is_memsize_b(ex_d_is_memsize_b),
    .ex_d_is_memsize_bu(ex_d_is_memsize_bu),
    .ex_d_is_memsize_h(ex_d_is_memsize_h),
    .ex_d_is_memsize_hu(ex_d_is_memsize_hu),
    .ex_d_is_memsize_w(ex_d_is_memsize_w),
    .ex_d_branch_predict(ex_d_branch_predict),
    .ex_d_pht_idx(ex_d_pht_idx),
    .ex_d_jump_taken(ex_d_jump_taken),
    .ex_d_jaddr(ex_d_jaddr),
    .ex_d_trap_valid(ex_d_trap_valid),
    .ex_d_trap_mcause(ex_d_trap_mcause),
    .ex_d_trap_pc(ex_d_trap_pc),
    .ex_d_insn(ex_d_insn),
    .ex_d_intr(ex_d_intr),
    .ex_d_next_pc(ex_d_next_pc),
    .ex_d_csr_rdata(ex_d_csr_rdata),
    .ex_d_rs1_addr(ex_d_rs1_addr),
    .ex_d_rs2_addr(ex_d_rs2_addr),
    .ex_d_rs1_rdata(ex_d_rs1_rdata),
    .ex_d_rs2_rdata(ex_d_rs2_rdata),
    .ex_d_trap_insn(ex_d_trap_insn),
    .ex_d_trap_next_pc(ex_d_trap_next_pc),
    .ex_d_trap_rs1_addr(ex_d_trap_rs1_addr),
    .ex_d_trap_rs2_addr(ex_d_trap_rs2_addr),
    .ex_d_trap_rd_addr(ex_d_trap_rd_addr),
    .ex_d_trap_rs1_rdata(ex_d_trap_rs1_rdata),
    .ex_d_trap_rs2_rdata(ex_d_trap_rs2_rdata),
    .ex_d_trap_rd_wdata(ex_d_trap_rd_wdata),
    .mem_q_insn(mem_q_insn),
    .mem_q_intr(mem_q_intr),
    .mem_q_next_pc(mem_q_next_pc),
    .mem_q_csr_rdata(mem_q_csr_rdata),
    .mem_q_rs1_addr(mem_q_rs1_addr),
    .mem_q_rs2_addr(mem_q_rs2_addr),
    .mem_q_rs1_rdata(mem_q_rs1_rdata),
    .mem_q_rs2_rdata(mem_q_rs2_rdata),
    .mem_q_trap_insn(mem_q_trap_insn),
    .mem_q_trap_next_pc(mem_q_trap_next_pc),
    .mem_q_trap_rs1_addr(mem_q_trap_rs1_addr),
    .mem_q_trap_rs2_addr(mem_q_trap_rs2_addr),
    .mem_q_trap_rd_addr(mem_q_trap_rd_addr),
    .mem_q_trap_rs1_rdata(mem_q_trap_rs1_rdata),
    .mem_q_trap_rs2_rdata(mem_q_trap_rs2_rdata),
    .mem_q_trap_rd_wdata(mem_q_trap_rd_wdata),
    .mem_q_valid(mem_q_valid),
    .mem_q_pc(mem_q_pc),
    .mem_q_pc_plus_4(mem_q_pc_plus_4),
    .mem_q_rd_addr(mem_q_rd_addr),
    .mem_q_csr_addr(mem_q_csr_addr),
    .mem_q_csr_wdata(mem_q_csr_wdata),
    .mem_q_store_wdata(mem_q_store_wdata),
    .mem_q_alu_csr_result(mem_q_alu_csr_result),
    .mem_q_is_branch(mem_q_is_branch),
    .mem_q_is_jump(mem_q_is_jump),
    .mem_q_is_csr_write(mem_q_is_csr_write),
    .mem_q_is_csr_read(mem_q_is_csr_read),
    .mem_q_is_rd_write(mem_q_is_rd_write),
    .mem_q_is_mem_write(mem_q_is_mem_write),
    .mem_q_is_mem_read(mem_q_is_mem_read),
    .mem_q_is_jal(mem_q_is_jal),
    .mem_q_is_jalr(mem_q_is_jalr),
    .mem_q_is_memsize_b(mem_q_is_memsize_b),
    .mem_q_is_memsize_bu(mem_q_is_memsize_bu),
    .mem_q_is_memsize_h(mem_q_is_memsize_h),
    .mem_q_is_memsize_hu(mem_q_is_memsize_hu),
    .mem_q_is_memsize_w(mem_q_is_memsize_w),
    .mem_q_branch_predict(mem_q_branch_predict),
    .mem_q_pht_idx(mem_q_pht_idx),
    .mem_q_jump_taken(mem_q_jump_taken),
    .mem_q_jaddr(mem_q_jaddr),
    .mem_q_trap_valid(mem_q_trap_valid),
    .mem_q_trap_mcause(mem_q_trap_mcause),
    .mem_q_trap_pc(mem_q_trap_pc)
  );

//-------------------------------
// MEM/WB pipeline
//-------------------------------
  mem_wb_pipeline  mem_wb_pipeline_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .mem_wb_flush(mem_wb_flush),
    .mem_wb_stall(mem_wb_stall),
    .ex_mem_stall(ex_mem_stall),
    .mem_d_valid(mem_d_valid),
    .mem_d_rd_addr(mem_d_rd_addr),
    .mem_d_csr_addr(mem_d_csr_addr),
    .mem_d_csr_wdata(mem_d_csr_wdata),
    .mem_d_rd_wdata(mem_d_rd_wdata),
    .mem_d_pc_plus_4(mem_d_pc_plus_4),
    .mem_d_is_csr_write(mem_d_is_csr_write),
    .mem_d_is_csr_read(mem_d_is_csr_read),
    .mem_d_is_rd_write(mem_d_is_rd_write),
    .mem_d_trap_valid(mem_d_trap_valid),
    .mem_d_trap_mcause(mem_d_trap_mcause),
    .mem_d_trap_pc(mem_d_trap_pc),
    .mem_d_pc(mem_d_pc),
    .mem_d_next_pc(mem_d_next_pc),
    .mem_d_insn(mem_d_insn),
    .mem_d_intr(mem_d_intr),
    .mem_d_csr_rdata(mem_d_csr_rdata),
    .mem_d_mem_addr(mem_d_mem_addr),
    .mem_d_load_rdata(mem_d_load_rdata),
    .mem_d_rs1_addr(mem_d_rs1_addr),
    .mem_d_rs2_addr(mem_d_rs2_addr),
    .mem_d_rs1_rdata(mem_d_rs1_rdata),
    .mem_d_rs2_rdata(mem_d_rs2_rdata),
    .mem_d_load_rmask(mem_d_load_rmask),
    .mem_d_store_wmask(mem_d_store_wmask),
    .mem_d_store_wdata(mem_d_store_wdata),
    .mem_d_trap_insn(mem_d_trap_insn),
    .mem_d_trap_next_pc(mem_d_trap_next_pc),
    .mem_d_trap_rs1_addr(mem_d_trap_rs1_addr),
    .mem_d_trap_rs2_addr(mem_d_trap_rs2_addr),
    .mem_d_trap_rd_addr(mem_d_trap_rd_addr),
    .mem_d_trap_rs1_rdata(mem_d_trap_rs1_rdata),
    .mem_d_trap_rs2_rdata(mem_d_trap_rs2_rdata),
    .mem_d_trap_rd_wdata(mem_d_trap_rd_wdata),
    .wb_q_pc(wb_q_pc),
    .wb_q_next_pc(wb_q_next_pc),
    .wb_q_insn(wb_q_insn),
    .wb_q_intr(wb_q_intr),
    .wb_q_csr_rdata(wb_q_csr_rdata),
    .wb_q_mem_addr(wb_q_mem_addr),
    .wb_q_load_rdata(wb_q_load_rdata),
    .wb_q_rs1_addr(wb_q_rs1_addr),
    .wb_q_rs2_addr(wb_q_rs2_addr),
    .wb_q_rs1_rdata(wb_q_rs1_rdata),
    .wb_q_rs2_rdata(wb_q_rs2_rdata),
    .wb_q_load_rmask(wb_q_load_rmask),
    .wb_q_store_wmask(wb_q_store_wmask),
    .wb_q_store_wdata(wb_q_store_wdata),
    .wb_q_trap_insn(wb_q_trap_insn),
    .wb_q_trap_next_pc(wb_q_trap_next_pc),
    .wb_q_trap_rs1_addr(wb_q_trap_rs1_addr),
    .wb_q_trap_rs2_addr(wb_q_trap_rs2_addr),
    .wb_q_trap_rd_addr(wb_q_trap_rd_addr),
    .wb_q_trap_rs1_rdata(wb_q_trap_rs1_rdata),
    .wb_q_trap_rs2_rdata(wb_q_trap_rs2_rdata),
    .wb_q_trap_rd_wdata(wb_q_trap_rd_wdata),
    .wb_q_valid(wb_q_valid),
    .wb_q_rd_addr(wb_q_rd_addr),
    .wb_q_csr_addr(wb_q_csr_addr),
    .wb_q_csr_wdata(wb_q_csr_wdata),
    .wb_q_rd_wdata(wb_q_rd_wdata),
    .wb_q_pc_plus_4(wb_q_pc_plus_4),
    .wb_q_is_csr_write(wb_q_is_csr_write),
    .wb_q_is_csr_read(wb_q_is_csr_read),
    .wb_q_is_rd_write(wb_q_is_rd_write),
    .wb_q_trap_valid(wb_q_trap_valid),
    .wb_q_trap_mcause(wb_q_trap_mcause),
    .wb_q_trap_pc(wb_q_trap_pc)
  );



  //*****************************************************************
  //
  //
  // REGISTER FILE
  //
  //
  //*****************************************************************

 riscv_regfile  riscv_regfile_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .id_rs1_addr(id_rs1_addr),
    .id_rs2_addr(id_rs2_addr),
    .wb_q_is_rd_write(wb_q_is_rd_write),
    .wb_rd_addr(wb_rd_addr),
    .wb_rd_wdata(wb_rd_wdata),
    .regfile_rs1_rdata(regfile_rs1_rdata),
    .regfile_rs2_rdata(regfile_rs2_rdata)
  );

  //*****************************************************************
  //
  //
  // CSR FILE
  //
  //
  //*****************************************************************
  csr_file csr_file_inst (
    .clk_i            (clk_i            ),
    .rst_i            (rst_i            ),
    .id_csr_addr      (id_csr_addr      ),
    .csrfile_rdata    (csrfile_rdata    ),
    .wb_q_valid       (wb_q_valid       ),
    .wb_q_trap_valid  (wb_q_trap_valid  ),
    .wb_q_is_csr_write(wb_q_is_csr_write),
    .wb_q_is_csr_read (wb_q_is_csr_read ),
    .wb_csr_addr      (wb_csr_addr      ),
    .wb_csr_wdata     (wb_csr_wdata     ),
    .wb_trap_pc       (wb_trap_pc       ),
    .wb_trap_mcause   (wb_trap_mcause   ),
    .ex_q_valid       (ex_q_valid       ),
    .mem_q_valid      (mem_q_valid      ),
    .wb_csr_rmask           (wb_csr_rmask           ),
    .wb_csr_wmask     (wb_csr_wmask     ),
    .trap_handler_addr(trap_handler_addr)
  );



  //*****************************************************************
  //
  //
  // HAZARD UNIT
  //
  //
  //*****************************************************************
  hazard_ctrl hazard_ctrl_inst (
    .id_rs1_addr          (id_rs1_addr          ),
    .id_rs2_addr          (id_rs2_addr          ),
    .ex_q_rs1_addr        (ex_q_rs1_addr        ),
    .ex_q_rs2_addr        (ex_q_rs2_addr        ),
    .ex_q_rd_addr         (ex_q_rd_addr         ),
    .mem_q_rd_addr        (mem_q_rd_addr        ),
    .wb_q_rd_addr         (wb_q_rd_addr         ),
    .ex_q_is_mem_read     (ex_q_is_mem_read     ),
    .mem_q_is_rd_write    (mem_q_is_rd_write    ),
    .wb_q_is_rd_write     (wb_q_is_rd_write     ),
    .mem_q_jump_taken     (mem_q_jump_taken     ),
    .mem_q_is_branch      (mem_q_is_branch      ),
    .mem_branch_mispredict(mem_branch_mispredict),
    .id_predict_btaken    (id_predict_btaken    ),
    .ex_q_trap_valid      (ex_q_trap_valid      ),
    .mem_q_trap_valid     (mem_q_trap_valid     ),
    .wb_q_trap_valid      (wb_q_trap_valid      ),
    .dmem_periph_req      (dmem_periph_req      ),
    .mem_done_i           (mem_done_i           ),
    .if_id_stall          (if_id_stall          ),
    .id_ex_stall          (id_ex_stall          ),
    .ex_mem_stall         (ex_mem_stall         ),
    .mem_wb_stall         (mem_wb_stall         ),
    .if_id_flush          (if_id_flush          ),
    .id_ex_flush          (id_ex_flush          ),
    .ex_mem_flush         (ex_mem_flush         ),
    .mem_wb_flush         (mem_wb_flush         ),
    .id_forward_rs1       (id_forward_rs1       ),
    .id_forward_rs2       (id_forward_rs2       ),
    .ex_forward_rs1_sel   (ex_forward_rs1_sel   ),
    .ex_forward_rs2_sel   (ex_forward_rs2_sel   )
  );

  //*****************************************************************
  //
  //
  // FORMAL VERIFICATION
  //
  //
  //*****************************************************************

`ifdef RISCV_FORMAL

riscv_formal_if  riscv_formal_if_inst (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .mem_wb_stall(mem_wb_stall),
    .trap_handler_addr(trap_handler_addr),
    .wb_csr_wmask(wb_csr_wmask),
    .wb_csr_rmask(wb_csr_rmask),
    .wb_q_pc(wb_q_pc),
    .wb_q_next_pc(wb_q_next_pc),
    .wb_q_insn(wb_q_insn),
    .wb_q_valid(wb_q_valid),
    .wb_q_trap_valid(wb_q_trap_valid),
    .wb_q_intr(wb_q_intr),
    .wb_q_rs1_addr(wb_q_rs1_addr),
    .wb_q_rs2_addr(wb_q_rs2_addr),
    .wb_q_rs1_rdata(wb_q_rs1_rdata),
    .wb_q_rs2_rdata(wb_q_rs2_rdata),
    .wb_q_is_rd_write(wb_q_is_rd_write),
    .wb_rd_addr(wb_rd_addr),
    .wb_rd_wdata(wb_rd_wdata),
    .wb_csr_addr(wb_csr_addr),
    .wb_q_csr_rdata(wb_q_csr_rdata),
    .wb_q_csr_wdata(wb_q_csr_wdata),
    .wb_q_is_csr_read(wb_q_is_csr_read),
    .wb_q_is_csr_write(wb_q_is_csr_write),
    .wb_q_mem_addr(wb_q_mem_addr),
    .wb_q_load_rdata(wb_q_load_rdata),
    .wb_q_store_wdata(wb_q_store_wdata),
    .wb_q_load_rmask(wb_q_load_rmask),
    .wb_q_store_wmask(wb_q_store_wmask),
    .wb_q_trap_insn(wb_q_trap_insn),
    .wb_q_trap_pc(wb_q_trap_pc),
    .wb_q_trap_next_pc(wb_q_trap_next_pc),
    .wb_q_trap_rs1_addr(wb_q_trap_rs1_addr),
    .wb_q_trap_rs2_addr(wb_q_trap_rs2_addr),
    .wb_q_trap_rd_addr(wb_q_trap_rd_addr),
    .wb_q_trap_rs1_rdata(wb_q_trap_rs1_rdata),
    .wb_q_trap_rs2_rdata(wb_q_trap_rs2_rdata),
    .wb_q_trap_rd_wdata(wb_q_trap_rd_wdata),
    .rvfi_valid(rvfi_valid),
    .rvfi_order(rvfi_order),
    .rvfi_insn(rvfi_insn),
    .rvfi_trap(rvfi_trap),
    .rvfi_halt(rvfi_halt),
    .rvfi_intr(rvfi_intr),
    .rvfi_mode(rvfi_mode),
    .rvfi_ixl(rvfi_ixl),
    .rvfi_rs1_addr(rvfi_rs1_addr),
    .rvfi_rs2_addr(rvfi_rs2_addr),
    .rvfi_rs1_rdata(rvfi_rs1_rdata),
    .rvfi_rs2_rdata(rvfi_rs2_rdata),
    .rvfi_rd_addr(rvfi_rd_addr),
    .rvfi_rd_wdata(rvfi_rd_wdata),
    .rvfi_pc_rdata(rvfi_pc_rdata),
    .rvfi_pc_wdata(rvfi_pc_wdata),
    .rvfi_mem_addr(rvfi_mem_addr),
    .rvfi_mem_rdata(rvfi_mem_rdata),
    .rvfi_mem_wdata(rvfi_mem_wdata),
    .rvfi_mem_rmask(rvfi_mem_rmask),
    .rvfi_mem_wmask(rvfi_mem_wmask),
    .rvfi_csr_mcycle_rdata(rvfi_csr_mcycle_rdata),
    .rvfi_csr_mcycle_wdata(rvfi_csr_mcycle_wdata),
    .rvfi_csr_mcycle_rmask(rvfi_csr_mcycle_rmask),
    .rvfi_csr_mcycle_wmask(rvfi_csr_mcycle_wmask),
    .rvfi_csr_minstret_rdata(rvfi_csr_minstret_rdata),
    .rvfi_csr_minstret_wdata(rvfi_csr_minstret_wdata),
    .rvfi_csr_minstret_rmask(rvfi_csr_minstret_rmask),
    .rvfi_csr_minstret_wmask(rvfi_csr_minstret_wmask),
    .rvfi_csr_mcause_rdata(rvfi_csr_mcause_rdata),
    .rvfi_csr_mcause_wdata(rvfi_csr_mcause_wdata),
    .rvfi_csr_mcause_rmask(rvfi_csr_mcause_rmask),
    .rvfi_csr_mcause_wmask(rvfi_csr_mcause_wmask),
    .rvfi_csr_mtvec_rdata(rvfi_csr_mtvec_rdata),
    .rvfi_csr_mtvec_wdata(rvfi_csr_mtvec_wdata),
    .rvfi_csr_mtvec_rmask(rvfi_csr_mtvec_rmask),
    .rvfi_csr_mtvec_wmask(rvfi_csr_mtvec_wmask),
    .rvfi_csr_mepc_rdata(rvfi_csr_mepc_rdata),
    .rvfi_csr_mepc_wdata(rvfi_csr_mepc_wdata),
    .rvfi_csr_mepc_rmask(rvfi_csr_mepc_rmask),
    .rvfi_csr_mepc_wmask(rvfi_csr_mepc_wmask)
  );
`endif


endmodule
